* Extracted by KLayout with SKY130 LVS runset on : 02/09/2023 21:00

.SUBCKT uldp
X$1 VN VP \$I1 VP VP VP VP VP MOSFET
X$2 VP Contact$2
X$3 VP Contact$1
X$4 VP \$I1 VN VN VN VN VN VN sky130_gnd MOSFET$1
X$5 VN Contact
X$6 VN Contact$1
.ENDS uldp

.SUBCKT Contact$2 \$1
.ENDS Contact$2

.SUBCKT Contact \$1
.ENDS Contact

.SUBCKT Contact$1 \$1
.ENDS Contact$1

.SUBCKT MOSFET$1 \$1 \$2 \$3 \$4 \$5 \$6 \$7 \$8 sky130_gnd
M$1 \$3 \$1 \$2 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1.5 AS=0.42
+ AD=0.2025 PS=3.56 PD=1.77
M$2 \$2 \$1 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1.5 AS=0.2025
+ AD=0.2025 PS=1.77 PD=1.77
M$3 \$4 \$1 \$2 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1.5 AS=0.2025
+ AD=0.2025 PS=1.77 PD=1.77
M$4 \$2 \$1 \$5 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1.5 AS=0.2025
+ AD=0.2025 PS=1.77 PD=1.77
M$5 \$5 \$1 \$2 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1.5 AS=0.2025
+ AD=0.2025 PS=1.77 PD=1.77
M$6 \$2 \$1 \$6 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1.5 AS=0.2025
+ AD=0.2025 PS=1.77 PD=1.77
M$7 \$6 \$1 \$2 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1.5 AS=0.2025
+ AD=0.2025 PS=1.77 PD=1.77
M$8 \$2 \$1 \$7 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1.5 AS=0.2025
+ AD=0.2025 PS=1.77 PD=1.77
M$9 \$7 \$1 \$2 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1.5 AS=0.2025
+ AD=0.2025 PS=1.77 PD=1.77
M$10 \$2 \$1 \$8 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1.5 AS=0.2025
+ AD=0.42 PS=1.77 PD=3.56
.ENDS MOSFET$1

.SUBCKT MOSFET \$1 \$2 \$3 \$4 \$5 \$6 \$7 \$8
M$1 \$2 \$1 \$3 \$9 sky130_fd_pr__pfet_01v8_lvt L=0.5 W=2 AS=0.56 AD=0.27
+ PS=4.56 PD=2.27
M$2 \$3 \$1 \$4 \$9 sky130_fd_pr__pfet_01v8_lvt L=0.5 W=2 AS=0.27 AD=0.27
+ PS=2.27 PD=2.27
M$3 \$4 \$1 \$3 \$9 sky130_fd_pr__pfet_01v8_lvt L=0.5 W=2 AS=0.27 AD=0.27
+ PS=2.27 PD=2.27
M$4 \$3 \$1 \$5 \$9 sky130_fd_pr__pfet_01v8_lvt L=0.5 W=2 AS=0.27 AD=0.27
+ PS=2.27 PD=2.27
M$5 \$5 \$1 \$3 \$9 sky130_fd_pr__pfet_01v8_lvt L=0.5 W=2 AS=0.27 AD=0.27
+ PS=2.27 PD=2.27
M$6 \$3 \$1 \$6 \$9 sky130_fd_pr__pfet_01v8_lvt L=0.5 W=2 AS=0.27 AD=0.27
+ PS=2.27 PD=2.27
M$7 \$6 \$1 \$3 \$9 sky130_fd_pr__pfet_01v8_lvt L=0.5 W=2 AS=0.27 AD=0.27
+ PS=2.27 PD=2.27
M$8 \$3 \$1 \$7 \$9 sky130_fd_pr__pfet_01v8_lvt L=0.5 W=2 AS=0.27 AD=0.27
+ PS=2.27 PD=2.27
M$9 \$7 \$1 \$3 \$9 sky130_fd_pr__pfet_01v8_lvt L=0.5 W=2 AS=0.27 AD=0.27
+ PS=2.27 PD=2.27
M$10 \$3 \$1 \$8 \$9 sky130_fd_pr__pfet_01v8_lvt L=0.5 W=2 AS=0.27 AD=0.56
+ PS=2.27 PD=4.56
.ENDS MOSFET
